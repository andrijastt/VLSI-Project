module deb;

endmodule
