module ps2;

endmodule
