module hex;

endmodule
